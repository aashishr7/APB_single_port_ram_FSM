package ram_env_pkg;

`include "seq_item.sv"
`include "uvm_sequence.sv"
`include "uvm_sequencer.sv"
`include "uvm_driver.sv"
`include "uvm_monitor.sv"
`include "uvm_scb.sv"
`include "uvm_agent.sv"
`include "uvm_env.sv"

endpackage